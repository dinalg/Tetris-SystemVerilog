module font_rom ( input [6:0] addr,
						output [3:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        4'b0000, // 0
        4'b0000, // 1
        4'b0000, // 2
        4'b0000, // 3
         // code x01
        4'b0000, // 0 
        4'b0000, // 1  **
        4'b0110, // 2  **
        4'b0110, // 3    
         // code x02
        4'b0000, // 0 
        4'b0000, // 1 **
        4'b1100, // 2  **
        4'b0110, // 3    
         // code x03
        4'b0000, // 0 
        4'b0000, // 1 ****
        4'b0000, // 2 
        4'b1111, // 3    
         // code x04
        4'b0000, // 0 
        4'b0000, // 1   **
        4'b0011, // 2  **
        4'b0110, // 3 
         // code x05
        4'b0000, // 0 
        4'b0000, // 1   ***
        4'b0111, // 2     *
        4'b0001, // 3
         // code x06
        4'b0000, // 0 
        4'b0000, // 1  ***
        4'b1110, // 2  *
        4'b1000, // 3
         // code x07
        4'b0000, // 0 
        4'b0000, // 1 ***
        4'b1110, // 2  * 
        4'b0100, // 3  
         // code x08
        4'b0100, // 0 *
        4'b0100, // 1 *
        4'b0100, // 2 * 
        4'b0100, // 3 *
         // code x09
        4'b0000, // 0 	
        4'b0010, // 1  *
        4'b0110, // 2 ** 
        4'b0100, // 3 *
         // code x0a
        4'b0000, // 0 	
        4'b0100, // 1 *
        4'b0110, // 2 ** 
        4'b0010, // 3  *
         // code x0b
        4'b0000, // 0 	
        4'b0010, // 1  *
        4'b0010, // 2  * 
        4'b0110, // 3 **
         // code x0c
        4'b0000, // 0 	
        4'b0000, // 1 *
        4'b1000, // 2 *** 
        4'b1110, // 3   
         // code x0d
        4'b0000, // 0 	
        4'b1100, // 1 **
        4'b1000, // 2 * 
        4'b1000, // 3 *
         // code x0e
        4'b0000, // 0 	
        4'b0110, // 1 **
        4'b0010, // 2  * 
        4'b0010, // 3  *
        // code x0f
        4'b0000, // 0 	
        4'b0000, // 1   *
        4'b0010, // 2 *** 
        4'b1110, // 3  
         // code x10
        4'b0000, // 0 *	
        4'b0100, // 1 *
        4'b0100, // 2 ** 
        4'b0110, // 3
         // code x11
        4'b0000, // 0 	
        4'b0010, // 1  *
        4'b0110, // 2 ** 
        4'b0010, // 3  *
         // code x12
        4'b0000, // 0 	
        4'b0000, // 1  *
        4'b0100, // 2 *** 
        4'b1110, // 3     
         // code x13
        4'b0000, // 0 	
        4'b0100, // 1  *
        4'b0110, // 2  ** 
        4'b0100, // 3  *	
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  
		  4'b0000,
		  4'b0000,
		  4'b0000,
		  4'b0000,
//		  // code x14
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111111, // 2  *******
//        8'b11011011, // 3 ** ** **
//        8'b11011011, // 4 ** ** **
//        8'b11011011, // 5 ** ** **
//        8'b01111011, // 6  **** **
//        8'b00011011, // 7    ** **
//        8'b00011011, // 8    ** **
//        8'b00011011, // 9    ** **
//        8'b00011011, // a    ** **
//        8'b00011011, // b    ** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x15
//        8'b00000000, // 0
//        8'b01111100, // 1  *****
//        8'b11000110, // 2 **   **
//        8'b01100000, // 3  **
//        8'b00111000, // 4   ***
//        8'b01101100, // 5  ** **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b01101100, // 8  ** **
//        8'b00111000, // 9   ***
//        8'b00001100, // a     **
//        8'b11000110, // b **   **
//        8'b01111100, // c  *****
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x16
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b11111110, // 8 *******
//        8'b11111110, // 9 *******
//        8'b11111110, // a *******
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x17
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00111100, // 3   ****
//        8'b01111110, // 4  ******
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b01111110, // 8  ******
//        8'b00111100, // 9   ****
//        8'b00011000, // a    **
//        8'b01111110, // b  ******
//        8'b00110000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x18
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00111100, // 3   ****
//        8'b01111110, // 4  ******
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x19
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b01111110, // 9  ******
//        8'b00111100, // a   ****
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00011000, // 5    **
//        8'b00001100, // 6     **
//        8'b11111110, // 7 *******
//        8'b00001100, // 8     **
//        8'b00011000, // 9    **
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00110000, // 5   **
//        8'b01100000, // 6  **
//        8'b11111110, // 7 *******
//        8'b01100000, // 8  **
//        8'b00110000, // 9   **
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b11000000, // 6 **
//        8'b11000000, // 7 **
//        8'b11000000, // 8 **
//        8'b11111110, // 9 *******
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00100100, // 5   *  *
//        8'b01100110, // 6  **  **
//        8'b11111111, // 7 ********
//        8'b01100110, // 8  **  **
//        8'b00100100, // 9   *  *
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00010000, // 4    *
//        8'b00111000, // 5   ***
//        8'b00111000, // 6   ***
//        8'b01111100, // 7  *****
//        8'b01111100, // 8  *****
//        8'b11111110, // 9 *******
//        8'b11111110, // a *******
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x1f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b11111110, // 4 *******
//        8'b11111110, // 5 *******
//        8'b01111100, // 6  *****
//        8'b01111100, // 7  *****
//        8'b00111000, // 8   ***
//        8'b00111000, // 9   ***
//        8'b00010000, // a    *
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x20
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x21
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00111100, // 3   ****
//        8'b00111100, // 4   ****
//        8'b00111100, // 5   ****
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00000000, // 9
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x22
//        8'b00000000, // 0
//        8'b01100110, // 1  **  **
//        8'b01100110, // 2  **  **
//        8'b01100110, // 3  **  **
//        8'b00100100, // 4   *  *
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x23
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b01101100, // 3  ** **
//        8'b01101100, // 4  ** **
//        8'b11111110, // 5 *******
//        8'b01101100, // 6  ** **
//        8'b01101100, // 7  ** **
//        8'b01101100, // 8  ** **
//        8'b11111110, // 9 *******
//        8'b01101100, // a  ** **
//        8'b01101100, // b  ** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x24
//        8'b00011000, // 0     **
//        8'b00011000, // 1     **
//        8'b01111100, // 2   *****
//        8'b11000110, // 3  **   **
//        8'b11000010, // 4  **    *
//        8'b11000000, // 5  **
//        8'b01111100, // 6   *****
//        8'b00000110, // 7       **
//        8'b00000110, // 8       **
//        8'b10000110, // 9  *    **
//        8'b11000110, // a  **   **
//        8'b01111100, // b   *****
//        8'b00011000, // c     **
//        8'b00011000, // d     **
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x25
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b11000010, // 4 **    *
//        8'b11000110, // 5 **   **
//        8'b00001100, // 6     **
//        8'b00011000, // 7    **
//        8'b00110000, // 8   **
//        8'b01100000, // 9  **
//        8'b11000110, // a **   **
//        8'b10000110, // b *    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x26
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111000, // 2   ***
//        8'b01101100, // 3  ** **
//        8'b01101100, // 4  ** **
//        8'b00111000, // 5   ***
//        8'b01110110, // 6  *** **
//        8'b11011100, // 7 ** ***
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01110110, // b  *** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x27
//        8'b00000000, // 0
//        8'b00110000, // 1   **
//        8'b00110000, // 2   **
//        8'b00110000, // 3   **
//        8'b01100000, // 4  **
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x28
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00001100, // 2     **
//        8'b00011000, // 3    **
//        8'b00110000, // 4   **
//        8'b00110000, // 5   **
//        8'b00110000, // 6   **
//        8'b00110000, // 7   **
//        8'b00110000, // 8   **
//        8'b00110000, // 9   **
//        8'b00011000, // a    **
//        8'b00001100, // b     **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x29
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00110000, // 2   **
//        8'b00011000, // 3    **
//        8'b00001100, // 4     **
//        8'b00001100, // 5     **
//        8'b00001100, // 6     **
//        8'b00001100, // 7     **
//        8'b00001100, // 8     **
//        8'b00001100, // 9     **
//        8'b00011000, // a    **
//        8'b00110000, // b   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01100110, // 5  **  **
//        8'b00111100, // 6   ****
//        8'b11111111, // 7 ********
//        8'b00111100, // 8   ****
//        8'b01100110, // 9  **  **
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b01111110, // 7  ******
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00110000, // c   **
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b01111110, // 7  ******
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x2f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000010, // 4       *
//        8'b00000110, // 5      **
//        8'b00001100, // 6     **
//        8'b00011000, // 7    **
//        8'b00110000, // 8   **
//        8'b01100000, // 9  **
//        8'b11000000, // a **
//        8'b10000000, // b *
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x30
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11001110, // 5 **  ***
//        8'b11011110, // 6 ** ****
//        8'b11110110, // 7 **** **
//        8'b11100110, // 8 ***  **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x31
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2
//        8'b00111000, // 3
//        8'b01111000, // 4    **
//        8'b00011000, // 5   ***
//        8'b00011000, // 6  ****
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b01111110, // b    **
//        8'b00000000, // c    **
//        8'b00000000, // d  ******
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x32
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b00000110, // 4      **
//        8'b00001100, // 5     **
//        8'b00011000, // 6    **
//        8'b00110000, // 7   **
//        8'b01100000, // 8  **
//        8'b11000000, // 9 **
//        8'b11000110, // a **   **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x33
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b00000110, // 4      **
//        8'b00000110, // 5      **
//        8'b00111100, // 6   ****
//        8'b00000110, // 7      **
//        8'b00000110, // 8      **
//        8'b00000110, // 9      **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x34
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00001100, // 2     **
//        8'b00011100, // 3    ***
//        8'b00111100, // 4   ****
//        8'b01101100, // 5  ** **
//        8'b11001100, // 6 **  **
//        8'b11111110, // 7 *******
//        8'b00001100, // 8     **
//        8'b00001100, // 9     **
//        8'b00001100, // a     **
//        8'b00011110, // b    ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x35
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b11000000, // 3 **
//        8'b11000000, // 4 **
//        8'b11000000, // 5 **
//        8'b11111100, // 6 ******
//        8'b00000110, // 7      **
//        8'b00000110, // 8      **
//        8'b00000110, // 9      **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x36
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111000, // 2   ***
//        8'b01100000, // 3  **
//        8'b11000000, // 4 **
//        8'b11000000, // 5 **
//        8'b11111100, // 6 ******
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x37
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b11000110, // 3 **   **
//        8'b00000110, // 4      **
//        8'b00000110, // 5      **
//        8'b00001100, // 6     **
//        8'b00011000, // 7    **
//        8'b00110000, // 8   **
//        8'b00110000, // 9   **
//        8'b00110000, // a   **
//        8'b00110000, // b   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x38
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b01111100, // 6  *****
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x39
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b01111110, // 6  ******
//        8'b00000110, // 7      **
//        8'b00000110, // 8      **
//        8'b00000110, // 9      **
//        8'b00001100, // a     **
//        8'b01111000, // b  ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00110000, // b   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000110, // 3      **
//        8'b00001100, // 4     **
//        8'b00011000, // 5    **
//        8'b00110000, // 6   **
//        8'b01100000, // 7  **
//        8'b00110000, // 8   **
//        8'b00011000, // 9    **
//        8'b00001100, // a     **
//        8'b00000110, // b      **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111110, // 5  ******
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b01111110, // 8  ******
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b01100000, // 3  **
//        8'b00110000, // 4   **
//        8'b00011000, // 5    **
//        8'b00001100, // 6     **
//        8'b00000110, // 7      **
//        8'b00001100, // 8     **
//        8'b00011000, // 9    **
//        8'b00110000, // a   **
//        8'b01100000, // b  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x3f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b00001100, // 5     **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00000000, // 9
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x40
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11011110, // 6 ** ****
//        8'b11011110, // 7 ** ****
//        8'b11011110, // 8 ** ****
//        8'b11011100, // 9 ** ***
//        8'b11000000, // a **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x41
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00010000, // 2    *
//        8'b00111000, // 3   ***
//        8'b01101100, // 4  ** **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11111110, // 7 *******
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x42
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11111100, // b ******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x43
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b01100110, // 3  **  **
//        8'b11000010, // 4 **    *
//        8'b11000000, // 5 **
//        8'b11000000, // 6 **
//        8'b11000000, // 7 **
//        8'b11000000, // 8 **
//        8'b11000010, // 9 **    *
//        8'b01100110, // a  **  **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x44
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111000, // 2 *****
//        8'b01101100, // 3  ** **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01100110, // 6  **  **
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01101100, // a  ** **
//        8'b11111000, // b *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x45
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b01100110, // 3  **  **
//        8'b01100010, // 4  **   *
//        8'b01101000, // 5  ** *
//        8'b01111000, // 6  ****
//        8'b01101000, // 7  ** *
//        8'b01100000, // 8  **
//        8'b01100010, // 9  **   *
//        8'b01100110, // a  **  **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x46
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b01100110, // 3  **  **
//        8'b01100010, // 4  **   *
//        8'b01101000, // 5  ** *
//        8'b01111000, // 6  ****
//        8'b01101000, // 7  ** *
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x47
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b01100110, // 3  **  **
//        8'b11000010, // 4 **    *
//        8'b11000000, // 5 **
//        8'b11000000, // 6 **
//        8'b11011110, // 7 ** ****
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b01100110, // a  **  **
//        8'b00111010, // b   *** *
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x48
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11111110, // 6 *******
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x49
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011110, // 2    ****
//        8'b00001100, // 3     **
//        8'b00001100, // 4     **
//        8'b00001100, // 5     **
//        8'b00001100, // 6     **
//        8'b00001100, // 7     **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01111000, // b  ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11100110, // 2 ***  **
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01101100, // 5  ** **
//        8'b01111000, // 6  ****
//        8'b01111000, // 7  ****
//        8'b01101100, // 8  ** **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11110000, // 2 ****
//        8'b01100000, // 3  **
//        8'b01100000, // 4  **
//        8'b01100000, // 5  **
//        8'b01100000, // 6  **
//        8'b01100000, // 7  **
//        8'b01100000, // 8  **
//        8'b01100010, // 9  **   *
//        8'b01100110, // a  **  **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11100111, // 3 ***  ***
//        8'b11111111, // 4 ********
//        8'b11111111, // 5 ********
//        8'b11011011, // 6 ** ** **
//        8'b11000011, // 7 **    **
//        8'b11000011, // 8 **    **
//        8'b11000011, // 9 **    **
//        8'b11000011, // a **    **
//        8'b11000011, // b **    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11100110, // 3 ***  **
//        8'b11110110, // 4 **** **
//        8'b11111110, // 5 *******
//        8'b11011110, // 6 ** ****
//        8'b11001110, // 7 **  ***
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x50
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01100000, // 7  **
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x510
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11010110, // 9 ** * **
//        8'b11011110, // a ** ****
//        8'b01111100, // b  *****
//        8'b00001100, // c     **
//        8'b00001110, // d     ***
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x52
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01101100, // 7  ** **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x53
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b01100000, // 5  **
//        8'b00111000, // 6   ***
//        8'b00001100, // 7     **
//        8'b00000110, // 8      **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x54
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111111, // 2 ********
//        8'b11011011, // 3 ** ** **
//        8'b10011001, // 4 *  **  *
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x55
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x56
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11000011, // 7 **    **
//        8'b11000011, // 8 **    **
//        8'b01100110, // 9  **  **
//        8'b00111100, // a   ****
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x57
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11011011, // 7 ** ** **
//        8'b11011011, // 8 ** ** **
//        8'b11111111, // 9 ********
//        8'b01100110, // a  **  **
//        8'b01100110, // b  **  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//        
//         // code x58
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b01100110, // 4  **  **
//        8'b00111100, // 5   ****
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00111100, // 8   ****
//        8'b01100110, // 9  **  **
//        8'b11000011, // a **    **
//        8'b11000011, // b **    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x59
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b01100110, // 5  **  **
//        8'b00111100, // 6   ****
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111111, // 2 ********
//        8'b11000011, // 3 **    **
//        8'b10000110, // 4 *    **
//        8'b00001100, // 5     **
//        8'b00011000, // 6    **
//        8'b00110000, // 7   **
//        8'b01100000, // 8  **
//        8'b11000001, // 9 **     *
//        8'b11000011, // a **    **
//        8'b11111111, // b ********
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b00110000, // 3   **
//        8'b00110000, // 4   **
//        8'b00110000, // 5   **
//        8'b00110000, // 6   **
//        8'b00110000, // 7   **
//        8'b00110000, // 8   **
//        8'b00110000, // 9   **
//        8'b00110000, // a   **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b10000000, // 3 *
//        8'b11000000, // 4 **
//        8'b11100000, // 5 ***
//        8'b01110000, // 6  ***
//        8'b00111000, // 7   ***
//        8'b00011100, // 8    ***
//        8'b00001110, // 9     ***
//        8'b00000110, // a      **
//        8'b00000010, // b       *
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b00001100, // 3     **
//        8'b00001100, // 4     **
//        8'b00001100, // 5     **
//        8'b00001100, // 6     **
//        8'b00001100, // 7     **
//        8'b00001100, // 8     **
//        8'b00001100, // 9     **
//        8'b00001100, // a     **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5e
//        8'b00010000, // 0    *
//        8'b00111000, // 1   ***
//        8'b01101100, // 2  ** **
//        8'b11000110, // 3 **   **
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b11111111, // d ********
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x60
//        8'b00110000, // 0   **
//        8'b00110000, // 1   **
//        8'b00011000, // 2    **
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x61
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111000, // 5  ****
//        8'b00001100, // 6     **
//        8'b01111100, // 7  *****
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01110110, // b  *** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x62
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11100000, // 2  ***
//        8'b01100000, // 3   **
//        8'b01100000, // 4   **
//        8'b01111000, // 5   ****
//        8'b01101100, // 6   ** **
//        8'b01100110, // 7   **  **
//        8'b01100110, // 8   **  **
//        8'b01100110, // 9   **  **
//        8'b01100110, // a   **  **
//        8'b01111100, // b   *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x63
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111100, // 5  *****
//        8'b11000110, // 6 **   **
//        8'b11000000, // 7 **
//        8'b11000000, // 8 **
//        8'b11000000, // 9 **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x64
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011100, // 2    ***
//        8'b00001100, // 3     **
//        8'b00001100, // 4     **
//        8'b00111100, // 5   ****
//        8'b01101100, // 6  ** **
//        8'b11001100, // 7 **  **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01110110, // b  *** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x65
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111100, // 5  *****
//        8'b11000110, // 6 **   **
//        8'b11111110, // 7 *******
//        8'b11000000, // 8 **
//        8'b11000000, // 9 **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x66
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111000, // 2   ***
//        8'b01101100, // 3  ** **
//        8'b01100100, // 4  **  *
//        8'b01100000, // 5  **
//        8'b11110000, // 6 ****
//        8'b01100000, // 7  **
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x67
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01110110, // 5  *** **
//        8'b11001100, // 6 **  **
//        8'b11001100, // 7 **  **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01111100, // b  *****
//        8'b00001100, // c     **
//        8'b11001100, // d **  **
//        8'b01111000, // e  ****
//        8'b00000000, // f
//         // code x68
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11100000, // 2 ***
//        8'b01100000, // 3  **
//        8'b01100000, // 4  **
//        8'b01101100, // 5  ** **
//        8'b01110110, // 6  *** **
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x69
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00011000, // 3    **
//        8'b00000000, // 4
//        8'b00111000, // 5   ***
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x6a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000110, // 2      **
//        8'b00000110, // 3      **
//        8'b00000000, // 4
//        8'b00001110, // 5     ***
//        8'b00000110, // 6      **
//        8'b00000110, // 7      **
//        8'b00000110, // 8      **
//        8'b00000110, // 9      **
//        8'b00000110, // a      **
//        8'b00000110, // b      **
//        8'b01100110, // c  **  **
//        8'b01100110, // d  **  **
//        8'b00111100, // e   ****
//        8'b00000000, // f
//         // code x6b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11100000, // 2 ***
//        8'b01100000, // 3  **
//        8'b01100000, // 4  **
//        8'b01100110, // 5  **  **
//        8'b01101100, // 6  ** **
//        8'b01111000, // 7  ****
//        8'b01111000, // 8  ****
//        8'b01101100, // 9  ** **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x6c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111000, // 2   ***
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x6d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11100110, // 5 ***  **
//        8'b11111111, // 6 ********
//        8'b11011011, // 7 ** ** **
//        8'b11011011, // 8 ** ** **
//        8'b11011011, // 9 ** ** **
//        8'b11011011, // a ** ** **
//        8'b11011011, // b ** ** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x6e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11011100, // 5 ** ***
//        8'b01100110, // 6  **  **
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b01100110, // b  **  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x6f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111100, // 5  *****
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x70
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11011100, // 5 ** ***
//        8'b01100110, // 6  **  **
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b01111100, // b  *****
//        8'b01100000, // c  **
//        8'b01100000, // d  **
//        8'b11110000, // e ****
//        8'b00000000, // f
//         // code x71
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01110110, // 5  *** **
//        8'b11001100, // 6 **  **
//        8'b11001100, // 7 **  **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01111100, // b  *****
//        8'b00001100, // c     **
//        8'b00001100, // d     **
//        8'b00011110, // e    ****
//        8'b00000000, // f
//         // code x72
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11011100, // 5 ** ***
//        8'b01110110, // 6  *** **
//        8'b01100110, // 7  **  **
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x73
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b01111100, // 5  *****
//        8'b11000110, // 6 **   **
//        8'b01100000, // 7  **
//        8'b00111000, // 8   ***
//        8'b00001100, // 9     **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x74
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00010000, // 2    *
//        8'b00110000, // 3   **
//        8'b00110000, // 4   **
//        8'b11111100, // 5 ******
//        8'b00110000, // 6   **
//        8'b00110000, // 7   **
//        8'b00110000, // 8   **
//        8'b00110000, // 9   **
//        8'b00110110, // a   ** **
//        8'b00011100, // b    ***
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x75
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11001100, // 5 **  **
//        8'b11001100, // 6 **  **
//        8'b11001100, // 7 **  **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01110110, // b  *** **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x76
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11000011, // 7 **    **
//        8'b11000011, // 8 **    **
//        8'b01100110, // 9  **  **
//        8'b00111100, // a   ****
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x77
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11000011, // 7 **    **
//        8'b11011011, // 8 ** ** **
//        8'b11011011, // 9 ** ** **
//        8'b11111111, // a ********
//        8'b01100110, // b  **  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x78
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11000011, // 5 **    **
//        8'b01100110, // 6  **  **
//        8'b00111100, // 7   ****
//        8'b00011000, // 8    **
//        8'b00111100, // 9   ****
//        8'b01100110, // a  **  **
//        8'b11000011, // b **    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x79
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111110, // b  ******
//        8'b00000110, // c      **
//        8'b00001100, // d     **
//        8'b11111000, // e *****
//        8'b00000000, // f
//         // code x7a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00000000, // 4
//        8'b11111110, // 5 *******
//        8'b11001100, // 6 **  **
//        8'b00011000, // 7    **
//        8'b00110000, // 8   **
//        8'b01100000, // 9  **
//        8'b11000110, // a **   **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x7b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00001110, // 2     ***
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b01110000, // 6  ***
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00001110, // b     ***
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x7c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011000, // 2    **
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00000000, // 6
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x7d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01110000, // 2  ***
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00001110, // 6     ***
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b01110000, // b  ***
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x7e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01110110, // 2  *** **
//        8'b11011100, // 3 ** ***
//        8'b00000000, // 4
//        8'b00000000, // 5
//        8'b00000000, // 6
//        8'b00000000, // 7
//        8'b00000000, // 8
//        8'b00000000, // 9
//        8'b00000000, // a
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x7f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00000000, // 2
//        8'b00000000, // 3
//        8'b00010000, // 4    *
//        8'b00111000, // 5   ***
//        8'b01101100, // 6  ** **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11111110, // a *******
//        8'b00000000, // b
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000  // f
        };

	assign data = ROM[addr];

endmodule  